//Sync FIFO sequence library
package fifo_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"
     `include "fifo_defines.sv"
     `include "fifo_base_item.sv"
     `include "fifo_base_monitor.sv"
     `include "fifo_base_sequencer.sv"
     `include "fifo_virtual_sequencer.sv"
     `include "fifo_base_seq.sv"
     `include "fifo_virtual_seq.sv"
     `include "fifo_base_driver.sv"
     `include "fifo_base_agent.sv"
    // `include "fifo_scoreboard.sv"
     `include "fifo_base_env.sv"
     `include "fifo_base_test.sv"
     

endpackage : fifo_pkg