parameter int DATA_WIDTH=8;
parameter int MEM_SIZE=16;